-- For oppgave a)

library ieee;
use ieee.std_logic_1164.all;

entity delay_modified is 
    port (
        -- System Clock and Reset
        rst_n        : in  std_ulogic;
        mclk         : in  std_ulogic;
        indata       : in  std_ulogic_vector(7 downto 0);
        outdata      : out std_ulogic_vector(7 downto 0)
    );  
end delay_modified;

architecture rtl of delay_modified is 
    signal a, b, c: std_ulogic_vector(7 downto 0);

    -- we're gonna get a train of 'uu', unless we
    -- define initial values for the signals
    signal x1, x2: std_ulogic_vector(7 downto 0); 
begin  
    process (rst_n, mclk) is    
    begin
        -- if the reset line isn't held at cycle 0, then
        -- all signals *will* be unresolved and undefined
        if (rst_n = '0') then       
            a <= (others => '0');
            x1 <= (others => '0');
            b <= (others => '0');
            x2 <= (others => '0');
            c <= (others => '0');
        elsif rising_edge(mclk) then
            -- This is a "register process" with sequential "registers"
            -- that only change every rising edge, meaning that each
            -- "register" only "sees" the value of the preceding "register"
            -- from the previous clock cycle. In practical terms, this means
            -- that the value in 'indata' traverses each "register" every
            -- clock cycle.
            
            -- map 'a' to 'indata', reflecting an instantaneous change
            a  <= indata;

            -- map 'x1' to 'a'
            x1 <= a;

            -- map 'b' to 'x1'
            b  <= x1;

            -- map 'x2' to 'b'
            x2 <= b;

            -- map 'c' to 'x2'
            c  <= x2;
        end if;
    end process;

    -- (combinatorial logic)
    -- map 'outdata' to 'c', reflecting an instantaneous change
    outdata  <= c;
end rtl;
